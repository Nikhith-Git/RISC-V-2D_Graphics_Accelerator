module hlo();
endmodule

hlo test from mac pc
